cicsimgen tran

*Nothing here

.lib  "/home/mudasir/.volare/sky130B/libs.tech/ngspice/sky130.lib.spice" tt

.lib "../../../tech/ngspice/temperature.spi" Tt

.lib "../../../tech/ngspice/supply.spi" Vt


*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
.include ../../../work/xsch/RPLY_EX0.spice

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0     dc 0

IBP 0 IBPS_4U dc 4u 

V0 IBNS_20U 0 dc 1


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT IBPS_4U VSS IBNS_20U RPLY_EX0

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

.save v(IBPS_4U) v(VSS) v(IBNS_20U) i(V0)

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 100p 2n 0

tran 10p 10n 1p
write
quit

.endc

.end

