magic
tech sky130B
magscale 1 2
timestamp 1675615114
<< locali >>
rect -160 1478 -20 1662
rect 208 1482 348 1666
rect 1046 1480 1186 1664
rect 1418 1482 1558 1666
rect 2242 1480 2382 1664
rect 2614 1480 2754 1664
rect 3440 1482 3580 1666
rect 3814 1478 3954 1662
rect 4642 1480 4782 1664
rect 5014 1480 5154 1664
rect 6040 1480 6180 1664
rect 6414 1482 6554 1666
rect -80 1000 240 1040
rect 1140 1000 1460 1040
rect 2360 1000 2620 1040
rect 3540 1000 3800 1040
rect 4740 1000 5020 1040
rect 6120 1000 6460 1040
rect -300 900 6700 1000
<< metal1 >>
rect -6 2018 58 2020
rect 1680 2018 2080 2020
rect -6 1986 6402 2018
rect -7 1974 6402 1986
rect -6 1962 6402 1974
rect 1680 1960 2080 1962
rect 2480 1930 2520 1962
rect 3685 1885 3715 1930
rect 40 1580 140 1600
rect 40 1500 60 1580
rect 120 1500 140 1580
rect 1270 1560 1330 1566
rect 3670 1560 3730 1566
rect 1264 1500 1270 1560
rect 1330 1500 1336 1560
rect 40 1480 140 1500
rect 1270 1494 1330 1500
rect 3670 1494 3730 1500
rect 4870 1560 4930 1566
rect 4870 1494 4930 1500
rect 6270 1560 6330 1566
rect 6270 1494 6330 1500
rect 50 1161 130 1170
rect 180 1161 1210 1170
rect 1260 1161 1340 1170
rect 1390 1161 2410 1170
rect 2460 1161 2530 1170
rect 2590 1161 3600 1170
rect 3650 1161 3740 1170
rect 3790 1161 4810 1170
rect 4850 1161 4960 1170
rect 4980 1161 6210 1170
rect 6250 1161 6350 1170
rect 29 1149 6376 1161
rect 50 1140 130 1149
rect 180 1140 1210 1149
rect 1260 1140 1340 1149
rect 1390 1140 2410 1149
rect 2460 1140 2530 1149
rect 2590 1140 3600 1149
rect 3650 1140 3740 1149
rect 3790 1140 4810 1149
rect 4850 1140 4960 1149
rect 4980 1140 6210 1149
rect 6250 1140 6350 1149
<< via1 >>
rect 60 1500 120 1580
rect 1270 1500 1330 1560
rect 3670 1500 3730 1560
rect 4870 1500 4930 1560
rect 6270 1500 6330 1560
<< metal2 >>
rect 40 1580 140 1600
rect 40 1500 60 1580
rect 120 1560 140 1580
rect 1270 1560 1330 1566
rect 120 1500 1270 1560
rect 1330 1500 3670 1560
rect 3730 1500 4870 1560
rect 4930 1500 6270 1560
rect 6330 1500 6336 1560
rect 40 1480 140 1500
rect 1270 1494 1330 1500
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_0
timestamp 1674928262
transform 1 0 6297 0 1 1570
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_1
timestamp 1674928262
transform 1 0 90 0 1 1569
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_2
timestamp 1674928262
transform 1 0 1297 0 1 1570
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_3
timestamp 1674928262
transform 1 0 2497 0 1 1570
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_4
timestamp 1674928262
transform 1 0 3697 0 1 1570
box -297 -570 297 570
use sky130_fd_pr__nfet_01v8_5CE34N  sky130_fd_pr__nfet_01v8_5CE34N_5
timestamp 1674928262
transform 1 0 4897 0 1 1570
box -297 -570 297 570
<< labels >>
flabel metal1 -6 1962 1860 1980 0 FreeSans 288 0 0 0 IBPS_4U
port 1 nsew
flabel locali -300 900 6700 1000 0 FreeSans 288 0 0 0 VSS
port 2 nsew
flabel metal2 120 1500 1270 1560 0 FreeSans 288 0 0 0 IBNS_20U
port 3 nsew
<< end >>
